/**********************************************
______________                ______________
______________ \  /\  /|\  /| ______________
______________  \/  \/ | \/ | ______________
descript:
author : WM
Version: VERA.0.0
created: 2020-05-22 15:33:55 +0800
madified:
***********************************************/


package test_package;
parameter  NUM = 6;
//==========================================================================
//-------- define ----------------------------------------------------------
typedef struct {
logic [32-1:0]  op ;
logic [NUM-1:0]  pl ;
} s_ing;

typedef struct {
logic [32-1:0]  op ;
logic [NUM-1:0]  pl ;
} z_ing;

logic [32-1:0]  data ;
z_ing zing_v0;
s_ing s_ing_v1;

//==========================================================================
//-------- instance --------------------------------------------------------

//==========================================================================
//-------- expression ------------------------------------------------------
assign  zing_v0.op[9] = 0;

endpackage:test_package
