/**********************************************
_______________________________________ 
___________    Cook Darwin   __________    
_______________________________________
descript:
author : Cook.Darwin
Version: VERA.0.0
created: 2020-05-22 15:39:18 +0800
madified:
***********************************************/
`timescale 1ns/1ps

module test_struct#(
    parameter  NUM = 6
)();
//==========================================================================
//-------- define ----------------------------------------------------------
typedef union {
logic [32-1:0]  op ;
logic [NUM-1:0]  pl ;
} s_ing;

typedef struct packed{
logic [32-1:0]  op ;
logic [NUM-1:0]  pl ;
} z_ing;

z_ing zing_v0;
s_ing s_ing_v1;
z_ing zingx_v0 [9-1:0][32-1:0];

//==========================================================================
//-------- instance --------------------------------------------------------

//==========================================================================
//-------- expression ------------------------------------------------------

endmodule
