/**********************************************
_______________________________________ 
___________    Cook Darwin   __________    
_______________________________________
descript:
author : Cook.Darwin
Version: VERA.0.0
created: 2020-05-21 17:00:16 +0800
madified:
***********************************************/
`timescale 1ns/1ps

module test_foreach();
//==========================================================================
//-------- define ----------------------------------------------------------
logic [32-1:0]  data[32-1:0] ;

//==========================================================================
//-------- instance --------------------------------------------------------

//==========================================================================
//-------- expression ------------------------------------------------------
always_comb begin 
    foreach(data[i1])begin
        if(false)begin
             data[i1] = '0;
        end
        else begin
            foreach(data[i1][i2])begin
                 data[i1][i2] = '1;
            end
        end
    end
end

endmodule
