/**********************************************
______________                ______________
______________ \  /\  /|\  /| ______________
______________  \/  \/ | \/ | ______________
descript:
author : WM
Version: VERA.0.0
created: 2020-08-19 19:03:51 +0800
madified:
***********************************************/
`timescale 1ns/1ps

module a_test_md (
    input                   clock,
    input                   rst,
    axi_stream_inf.master   origin_inf
);

//==========================================================================
//-------- define ----------------------------------------------------------


//==========================================================================
//-------- instance --------------------------------------------------------

//==========================================================================
//-------- expression ------------------------------------------------------

endmodule
