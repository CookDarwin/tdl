/**********************************************
______________                ______________
______________ \  /\  /|\  /| ______________
______________  \/  \/ | \/ | ______________
descript:
author : WM
Version: VERA.0.0
created: 2020-08-19 14:57:59 +0800
madified:
***********************************************/
`timescale 1ns/1ps

module tb_test_top();
//==========================================================================
//-------- define ----------------------------------------------------------


//==========================================================================
//-------- instance --------------------------------------------------------
test_top rtl_top(
/* input clock */.sys_clock ( ),
/* output      */.odata     ( )
);
//==========================================================================
//-------- expression ------------------------------------------------------

endmodule
