/**********************************************
_______________________________________ 
___________    Cook Darwin   __________    
_______________________________________
descript:
author : Cook.Darwin
Version: VERA.0.0
created: 2020-08-19 15:56:21 +0800
madified:
***********************************************/
`timescale 1ns/1ps

module sdl_md (
    input                   clock,
    input                   rst_n,
    output logic[7:0]       odata,
    axi_stream_inf.slaver   asi_inf
);

//==========================================================================
//-------- define ----------------------------------------------------------


//==========================================================================
//-------- instance --------------------------------------------------------

//==========================================================================
//-------- expression ------------------------------------------------------

endmodule
