/**********************************************
______________                ______________
______________ \  /\  /|\  /| ______________
______________  \/  \/ | \/ | ______________
descript:
author : WM
Version: VERA.0.0
created: 2020-05-22 18:23:27 +0800
madified:
***********************************************/
`timescale 1ns/1ps
`include "define_macro.sv" 

module test_vcs_string#(
    `parameter_longstring(111) INIT_FILE = "ppppppppp"
)();
//==========================================================================
//-------- define ----------------------------------------------------------


//==========================================================================
//-------- instance --------------------------------------------------------

//==========================================================================
//-------- expression ------------------------------------------------------

endmodule
