/**********************************************
_______________________________________ 
___________    Cook Darwin   __________    
_______________________________________
descript:
author : Cook.Darwin
Version: VERA.0.0
created: xxxx.xx.xx
madified:
***********************************************/
`timescale 1ns/1ps

module exp_random #(
    parameter  PX = 67
)(
    output logic      param_random_b,
    output logic      int_random_b,
    output logic[9:0] rd_range
);

//==========================================================================
//-------- define ----------------------------------------------------------


//==========================================================================
//-------- instance --------------------------------------------------------

//==========================================================================
//-------- expression ------------------------------------------------------
initial begin
     param_random_b = ($urandom_range(0,99) <= PX);
     int_random_b = ($urandom_range(1,100) > 34);
     rd_range = $urandom_range(12,1000);
end

endmodule
