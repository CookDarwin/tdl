
module hdl_md #(
    parameter   DSIZE    =12
)(
    input                   clock,
    input                   rst_n,
    output logic[11:0]      odata,    
    axi_stream_inf.master   in_axis
);


endmodule

