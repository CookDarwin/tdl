/**********************************************
______________                ______________
______________ \  /\  /|\  /| ______________
______________  \/  \/ | \/ | ______________
descript:
author : WM
Version: VERA.0.0
created: 2020-08-19 10:31:59 +0800
madified:
***********************************************/


package head_package;
parameter  HDSIZE = 8;
//==========================================================================
//-------- define ----------------------------------------------------------
typedef struct {
logic [4-1:0]  idata ;
logic valid;
} s_head;


//==========================================================================
//-------- instance --------------------------------------------------------

//==========================================================================
//-------- expression ------------------------------------------------------

endpackage:head_package
