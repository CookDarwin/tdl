/**********************************************
______________                ______________
______________ \  /\  /|\  /| ______________
______________  \/  \/ | \/ | ______________
descript:
author : WM
Version: VERA.0.0
created: 2020-06-10 11:18:14 +0800
madified:
***********************************************/
`timescale 1ns/1ps

module test_initial_assert ();
//==========================================================================
//-------- define ----------------------------------------------------------
logic ppx;

//==========================================================================
//-------- instance --------------------------------------------------------

//==========================================================================
//-------- expression ------------------------------------------------------
initial begin 
    assert(9)else begin
         $error("iiiiiiiiiiiii");
         $stop;
    end
     ppx = 1'b0;
end

endmodule
