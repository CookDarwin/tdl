/**********************************************
_______________________________________ 
___________    Cook Darwin   __________    
_______________________________________
descript:
author : Cook.Darwin
Version: VERA.0.0
created: xxxx.xx.xx
madified:
***********************************************/
`timescale 1ns/1ps

module tb_test_top();
//==========================================================================
//-------- define ----------------------------------------------------------
logic gl_clk;
string test_unit_region;
logic [0-1:0]  unit_pass_u ;
logic [0-1:0]  unit_pass_d ;

//==========================================================================
//-------- instance --------------------------------------------------------
test_top rtl_top(
/* input clock */.global_sys_clk (gl_clk )
);
//==========================================================================
//-------- expression ------------------------------------------------------
initial begin
     forever begin #(33ns);gl_clk = ~gl_clk;end;
end

endmodule
